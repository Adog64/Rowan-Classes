module Lab1(HEX0, SW);
	input [7:0] SW;
	output [7:0] HEX0;
	assign HEX0 = SW;
endmodule